module orgatee ( a ,b ,y );

input a ;
wire a ;
input b ;
wire b ;
output y ;
wire y ;
assign y = a|b ;

endmodule
